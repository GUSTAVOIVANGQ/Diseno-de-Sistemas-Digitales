module escalera ( 
	a,
	b,
	a1,
	b1,
	c1,
	x1,
	x2,
	x3,
	x4,
	c
	) ;

input  a;
input  b;
input  a1;
input  b1;
input  c1;
inout  x1;
inout  x2;
inout  x3;
inout  x4;
inout  c;
